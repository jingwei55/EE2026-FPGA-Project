`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03.04.2022 16:44:12
// Design Name: 
// Module Name: Landmarks
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Landmarks(input CLOCK, input clk1k, input pbu, pbd, pbl, pbr, pbc, SW14, input [12:0] pixel_index, input [2:0] layer, input [31:0] x, y, output reg [15:0] oled_data);
    parameter [31:0] a = 4; 
    wire map, zoo, birdpark, bthill, esplanade, changi, sentosa, flyer, garden, merlion, def0, def1, def2, def3, def4, def5, def6, def7, def8;
    reg [4:0] state = 0;
    wire [15:0] landmark [4:0];
    
    reg[15:0] flyer_data[0:6143];
    reg[15:0] bthill_data[0:6143];reg[15:0] sentosa_data[0:6143];
    reg[15:0] changi_data[0:6143];reg[15:0] gardens_data[0:6143];
    reg[15:0] birdpark_data[0:6143];reg[15:0] merlion_data[0:6143];
    reg[15:0] zoo_data[0:6143];
    initial begin
    $readmemh("flyer.mem", flyer_data);
    $readmemh("merlion.mem", merlion_data);
    $readmemh("gardens.mem", gardens_data);
    $readmemh("sentosa.mem", sentosa_data);
    $readmemh("bthill.mem", bthill_data);
    $readmemh("changi.mem", changi_data);
    $readmemh("birdpark.mem", birdpark_data);
    $readmemh("zoo.mem", zoo_data);
    end
    
    assign map = (y==a && (x>= 45 && x<=53)) || (y==a+1 && (x>= 44 && x<=54)) || (y==a+2 && (x>= 41 && x<=55)) || (y==a+3 && (x>= 41 && x<=55)) || (y==a+4 && ((x>= 28 && x<=31)||(x>=39 && x<=57)))
                    || (y==a+5 && ((x>= 28 && x<=31)||(x>= 39 && x<=57))) || (y==a+6 && ((x>= 25 && x<=32)||(x>= 39 && x<=58))) || (y==a+7 && ((x>= 24 && x<=32)||(x>= 37 && x<=58))) || (y==a+8 && (x>= 23 && x<=57))
                    || (y==a+9 && ((x>= 21 && x<=57)||(x>=60 && x<=63))) 
                    || (y==a+10 && ((x>= 19 && x<=55)||(x>= 59 && x<=63)||(x>= 72 && x<=76))) 
                    || (y==a+11 && ((x>= 19 && x<=55)||(x>= 59 && x<=63)||(x==65)||(x>= 72 && x<=76))) 
                    || (y==a+12 && ((x>= 19 && x<=53)||(x>= 57 && x<=65)||(x>=67 && x<=68)||(x>= 73 && x<=81)))                
                    || (y==a+13 && ((x>= 19 && x<=51)||(x>= 56 && x<=65)||(x>=67 && x<=68)||(x>= 77 && x<=83))) 
                    || (y==a+14 && ((x>= 18 && x<=51)||(x>= 53 && x<=69)||(x>= 78 && x<=81)))
                    || (y==a+15 && ((x>= 18 && x<=49)||(x>= 53 && x<=69)||(x>= 78 && x<=81))) || (y==a+16 && (x>= 17 && x<=72)) || (y==a+17 && ((x>= 17 && x<=73)||(x>=83 && x<=85))) || (y==a+18 && ((x>= 17 && x<=73)||(x>=83 && x<=85))) 
                    || (y==a+19 && ((x>= 17 && x<=75)||(x>=82 && x<=89))) || (y==a+20 && ((x>= 16 && x<=77)||(x>=80 && x<=88))) || (y==a+21 && (x>= 16 && x<=89)) || (y==a+22 && (x>= 16 && x<=89)) || (y==a+23 && (x>= 13 && x<=88)) 
                    || (y==a+24 && (x>= 13 && x<=88)) || (y==a+25 && (x>= 12 && x<=89)) || (y==a+26 && (x>= 12 && x<=89)) || (y==a+27 && (x>= 11 && x<=89)) || (y==a+28 && (x>= 11 && x<=89)) || (y==a+29 && (x>= 11 && x<=89)) || (y==a+30 && (x>= 11 && x<=88)) || (y==a+31 && (x>= 10 && x<=88)) || (y==a+32 && (x>= 10 && x<=88)) || (y==a+33 && (x>= 10 && x<=87)) || (y==a+34 && (x>= 10 && x<=87)) || (y==a+35 && (x>= 10 && x<=90)) 
                    || (y==a+36 && (x>= 9 && x<=91)) || (y==a+37 && ((x>= 9 && x<=10)||(x>=13 && x<=77))) || (y==a+38 && ((x>= 9 && x<=10)||(x>=16 && x<=24)||(x>=30 && x<=71))) || (y==a+39 && ((x>= 8 && x<=11)||(x>=16 && x<=18)||(x>=34 && x<=67))) || (y==a+40 && ((x>= 8 && x<=11)||(x>=16 && x<=18)||(x>=34 && x<=67))) || (y==a+41 && ((x>= 8 && x<=12)||(x>=16 && x<=18)||(x>=27 && x<=29)||(x>=37 && x<=65))) || (y==a+42 && ((x>= 8 && x<=12)||(x>=24 && x<=29)||(x>=39 && x<=63))) 
                    || (y==a+43 && ((x>= 9 && x<=12)||(x>=24 && x<=30)||(x>=35 && x<=38)||(x>=40 && x<=60))) || (y==a+44 && ((x>= 9 && x<=12)||(x>=24 && x<=30)||(x>=35 && x<=38)||(x>=40 && x<=60))) || (y==a+45 && ((x>= 19 && x<=20)||(x>=23 && x<=33)||(x>=36 && x<=39)||(x>=42 && x<=59))) || (y==a+46 && ((x>= 18 && x<=21)||(x>=23 && x<=29)||(x==32)||(x>=37 && x<=39)||(x>=45 && x<=58))) || (y==a+47 && ((x>= 18 && x<=21)||(x>=23 && x<=29)||(x==32)||(x>=37 && x<=39)||(x>=45 && x<=58))) 
                    || (y==a+48 && ((x>= 17 && x<=26)||(x>=28 && x<=30)||(x>=46 && x<=54))) || (y==a+49 && ((x>= 16 && x<=24)||(x>=49 && x<=50))) || (y==a+50 && ((x>= 17 && x<=22)||(x>=24 && x<=26)||(x>=47 && x<=50)||(x>=52 && x<=54))) || (y==a+51 && ((x>= 17 && x<=21)||(x>=48 && x<=55))) || (y==a+52 && ((x>= 18 && x<=20)||(x>=51 && x<=54)))
                    || (y==a+53 && ((x>= 18 && x<=20)||(x>=51 && x<=54))) || (y==a+54 && ((x>= 18 && x<=20)||(x==52))) || (y==a+55 && ((x>= 18 && x<=20)||(x==52)));
                    
    assign merlion = (x == 61 && (y >= 41 - 1 && y <= 41 + 1)) || (y == 41 && (x== 61 - 1 || x== 61 + 1));
    assign flyer = (x == 67 && (y >= 42 - 1 && y <= 42 + 1)) || (y == 42 && (x== 67 - 1 || x== 67 + 1));
    assign garden = (x == 58 && (y >= 46 - 1 && y <= 46 + 1)) || (y == 46 && (x== 58 - 1 || x== 58 + 1));
    assign changi = (x == 84 && (y >= 31 - 1 && y <= 31 + 1)) || (y == 31 && (x== 84 - 1 || x== 84 + 1));
    assign bthill = (x == 46 && (y >= 32 - 1 && y <= 32 + 1)) || (y == 32 && (x== 46 - 1 || x== 46 + 1));
    assign sentosa = (x == 52 && (y >= 56 - 1 && y <= 56 + 1)) || (y == 56 && (x== 52 - 1 || x== 52 + 1));
    assign zoo = (x == 38 && (y >= 20 - 1 && y <= 20 + 1)) || (y == 20 && (x== 38 - 1 || x== 38 + 1));
    assign birdpark = (x == 25 && (y >= 37 - 1 && y <= 37 + 1)) || (y == 37 && (x== 25 - 1 || x== 25 + 1));   
    assign def0 =  merlion || flyer || garden || changi || bthill || sentosa || zoo || birdpark;
    assign def1 =  flyer || garden || changi || bthill || sentosa || zoo || birdpark;
    assign def2 =  merlion  || garden || changi || bthill || sentosa || zoo || birdpark;
    assign def3 =  merlion || flyer || changi || bthill || sentosa || zoo || birdpark;
    assign def4 =  merlion || flyer || garden || bthill || sentosa || zoo || birdpark;
    assign def5 =  merlion || flyer || garden || changi || sentosa || zoo || birdpark;
    assign def6 =  merlion || flyer || garden || changi || bthill || zoo || birdpark;
    assign def7 =  merlion || flyer || garden || changi || bthill || sentosa || birdpark;
    assign def8 =  merlion || flyer || garden || changi || bthill || sentosa || zoo;
    
    
    assign landmark[0] = map && ~def0;
    assign landmark[1] = map && ~def0; //merlion
    assign landmark[2] = map && ~def0; //flyer
    assign landmark[3] = map && ~def0; //garden
    assign landmark[4] = map && ~def0; //changi
    assign landmark[5] = map && ~def0; //bthill
    assign landmark[6] = map && ~def0; ///sentosa
    assign landmark[7] = map && ~def0; //zoo
    assign landmark[8] = map && ~def0; //birdpark
    
    assign landmark[9] = def0; //merlion photo here
    assign landmark[10] = def0; //flyer photo here
    assign landmark[11] = def0; //garden photo here
    assign landmark[12] = def0; //changi photo here
    assign landmark[13] = def0; //bthill photo here
    assign landmark[14] = def0; //sentosa photo here
    assign landmark[15] = def0; //zoo photo here
    assign landmark[16] = def0; //birdpark photo here
    
    always @ (posedge clk1k) begin
        if (SW14 && layer == 3) state <= 0; //reset
        else begin
        if (state == 0 && (pbu || pbr || pbc || pbl || pbd) && layer == 3)  state <= 5;
        else if (state == 5 && pbu && layer == 3) state <= 7; //bthill
        else if (state == 5 && pbd && layer == 3) state <= 3;
        else if (state == 5 && pbr && layer == 3) state <= 4;
        else if (state == 5 && pbl && layer == 3) state <= 8;
        else if (state == 5 && pbc && layer == 3) state <= 5+8;
        
        else if (state == 7 && pbd && layer == 3) state <= 5; //zoo
        else if (state == 7 && pbr && layer == 3) state <= 4;
        else if (state == 7 && pbl && layer == 3) state <= 8;
        else if (state == 7 && pbc && layer == 3) state <= 7+8;
        
        else if (state == 4 && pbu && layer == 3) state <= 7; //changi
        else if (state == 4 && pbd && layer == 3) state <= 2;
        else if (state == 4 && pbl && layer == 3) state <= 5;
        else if (state == 4 && pbc && layer == 3) state <= 4+8;
        
        else if (state == 2 && pbu && layer == 3) state <= 4; //flyer
        else if (state == 2 && pbr && layer == 3) state <= 4;
        else if (state == 2 && pbl && layer == 3) state <= 1;
        else if (state == 2 && pbc && layer == 3) state <= 2+8;
        
        else if (state == 3 && pbu && layer == 3) state <= 1; //garden
        else if (state == 3 && pbr && layer == 3) state <= 1;
        else if (state == 3 && pbl && layer == 3) state <= 8;
        else if (state == 3 && pbd && layer == 3) state <= 6;
        else if (state == 3 && pbc && layer == 3) state <= 3+8;
        
        else if (state == 6 && pbu && layer == 3) state <= 5; //sentosa
        else if (state == 6 && pbr && layer == 3) state <= 3;
        else if (state == 6 && pbl && layer == 3) state <= 8; 
        else if (state == 6 && pbc && layer == 3) state <= 6+8;
        
        else if (state == 8 && pbu && layer == 3) state <= 7; //birdpark
        else if (state == 8 && pbd && layer == 3) state <= 6;
        else if (state == 8 && pbr && layer == 3) state <= 5;
        else if (state == 8 && pbc && layer == 3) state <= 8+8;
        
        else if (state == 1 && pbu && layer == 3) state <= 5; //merlion
        else if (state == 1 && pbd && layer == 3) state <= 3;
        else if (state == 1 && pbr && layer == 3) state <= 2;
        else if (state == 1 && pbl && layer == 3) state <= 8;
        else if (state == 1 && pbc && layer == 3) state <= 1+8;
        
        else if (state >= 9 && state <= 16 && pbc && layer == 3) state <= 0; //return to default once picture is shown
        
        else state <= state;
        
        end
    end
    
    always @ (posedge CLOCK) begin
        if(state == 9)begin //merlion
            oled_data = merlion_data[pixel_index];
        end
                      
        else if(state == 10)begin
            oled_data = flyer_data[pixel_index];
        end
        
        else if(state == 11)begin
            oled_data = gardens_data[pixel_index];
        end
        
        else if(state ==12)begin
            oled_data = changi_data[pixel_index];
        end
        else if(state == 13)begin
            oled_data = bthill_data[pixel_index];        
        end
        else if(state == 14)begin
            oled_data = sentosa_data[pixel_index];
        end
        else if(state == 15) begin
            oled_data = zoo_data[pixel_index];
        end
        else if(state == 16)begin
            oled_data = birdpark_data[pixel_index];
        end
        else if(state >= 0 && state <= 8) begin
            oled_data = landmark[state] ? 16'b00000_111111_00000 : (state == 0 && def0) ? 16'b11111_000000_00000 
            : (state == 1 && def1) ? 16'b11111_000000_00000 : (state == 1 && merlion) ? 16'b11111_111111_00000 
            : (state == 2 && def2) ? 16'b11111_000000_00000 : (state == 2 && flyer) ? 16'b11111_111111_00000 
            : (state == 3 && def3) ? 16'b11111_000000_00000 : (state == 3 && garden) ? 16'b11111_111111_00000 
            : (state == 4 && def4) ? 16'b11111_000000_00000 : (state == 4 && changi) ? 16'b11111_111111_00000 
            : (state == 5 && def5) ? 16'b11111_000000_00000 : (state == 5 && bthill) ? 16'b11111_111111_00000 
            : (state == 6 && def6) ? 16'b11111_000000_00000 : (state == 6 && sentosa) ? 16'b11111_111111_00000 
            : (state == 7 && def7) ? 16'b11111_000000_00000 : (state == 7 && zoo) ? 16'b11111_111111_00000 
            : (state == 8 && def8) ? 16'b11111_000000_00000 : (state == 8 && birdpark) ? 16'b11111_111111_00000 : 0;
       end
    end
endmodule
