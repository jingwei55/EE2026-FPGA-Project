`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.04.2022 16:37:12
// Design Name: 
// Module Name: lockdown_animation
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module lockdown_animation(
    input CLOCK,
    input rst,
    input [12:0] pixel_index,
    output reg [15:0] oled_data
    );
    
always@(CLOCK)begin
    if (((pixel_index >= 0) && (pixel_index <= 2442)) || ((pixel_index >= 2444) && (pixel_index <= 2446)) || ((pixel_index >= 2450) && (pixel_index <= 2454)) || pixel_index == 2456 || ((pixel_index >= 2459) && (pixel_index <= 2529)) || ((pixel_index >= 2532) && (pixel_index <= 2537)) || pixel_index == 2539 || pixel_index == 2541 || pixel_index == 2543 || ((pixel_index >= 2545) && (pixel_index <= 2546)) || pixel_index == 2551 || ((pixel_index >= 2553) && (pixel_index <= 2554)) || ((pixel_index >= 2558) && (pixel_index <= 2614)) || ((pixel_index >= 2617) && (pixel_index <= 2624)) || pixel_index == 2627 || pixel_index == 2631 || pixel_index == 2634 || pixel_index == 2637 || pixel_index == 2639 || pixel_index == 2641 || pixel_index == 2643 || pixel_index == 2647 || pixel_index == 2649 || pixel_index == 2651 || ((pixel_index >= 2654) && (pixel_index <= 2708)) || ((pixel_index >= 2715) && (pixel_index <= 2721)) || pixel_index == 2723 || pixel_index == 2727 || pixel_index == 2732 || pixel_index == 2735 || pixel_index == 2737 || pixel_index == 2739 || pixel_index == 2743 || ((pixel_index >= 2750) && (pixel_index <= 2804)) || ((pixel_index >= 2806) && (pixel_index <= 2809)) || ((pixel_index >= 2811) && (pixel_index <= 2816)) || ((pixel_index >= 2829) && (pixel_index <= 2831)) || pixel_index == 2833 || ((pixel_index >= 2845) && (pixel_index <= 2900)) || ((pixel_index >= 2902) && (pixel_index <= 2905)) || ((pixel_index >= 2908) && (pixel_index <= 2988)) || ((pixel_index >= 2992) && (pixel_index <= 2996)) || ((pixel_index >= 3004) && (pixel_index <= 3006)) || ((pixel_index >= 3011) && (pixel_index <= 3013)) || ((pixel_index >= 3016) && (pixel_index <= 3017)) || pixel_index == 3021 || ((pixel_index >= 3026) && (pixel_index <= 3032)) || ((pixel_index >= 3036) && (pixel_index <= 3038)) || ((pixel_index >= 3041) && (pixel_index <= 3043)) || ((pixel_index >= 3046) && (pixel_index <= 3048)) || pixel_index == 3051 || ((pixel_index >= 3054) && (pixel_index <= 3056)) || ((pixel_index >= 3059) && (pixel_index <= 3084)) || ((pixel_index >= 3088) && (pixel_index <= 3092)) || ((pixel_index >= 3100) && (pixel_index <= 3101)) || ((pixel_index >= 3108) && (pixel_index <= 3109)) || pixel_index == 3112 || ((pixel_index >= 3116) && (pixel_index <= 3117)) || ((pixel_index >= 3124) && (pixel_index <= 3126)) || pixel_index == 3134 || ((pixel_index >= 3137) && (pixel_index <= 3139)) || ((pixel_index >= 3142) && (pixel_index <= 3143)) || pixel_index == 3147 || ((pixel_index >= 3151) && (pixel_index <= 3152)) || ((pixel_index >= 3155) && (pixel_index <= 3180)) || ((pixel_index >= 3184) && (pixel_index <= 3187)) || pixel_index == 3196 || ((pixel_index >= 3200) && (pixel_index <= 3202)) || ((pixel_index >= 3204) && (pixel_index <= 3205)) || ((pixel_index >= 3211) && (pixel_index <= 3213)) || ((pixel_index >= 3216) && (pixel_index <= 3217)) || pixel_index == 3221 || ((pixel_index >= 3225) && (pixel_index <= 3227)) || ((pixel_index >= 3230) && (pixel_index <= 3231)) || pixel_index == 3234 || pixel_index == 3239 || ((pixel_index >= 3242) && (pixel_index <= 3243)) || pixel_index == 3248 || ((pixel_index >= 3251) && (pixel_index <= 3276)) || ((pixel_index >= 3280) && (pixel_index <= 3283)) || pixel_index == 3292 || ((pixel_index >= 3295) && (pixel_index <= 3301)) || ((pixel_index >= 3306) && (pixel_index <= 3309)) || ((pixel_index >= 3312) && (pixel_index <= 3314)) || pixel_index == 3317 || ((pixel_index >= 3320) && (pixel_index <= 3323)) || pixel_index == 3327 || pixel_index == 3330 || pixel_index == 3335 || ((pixel_index >= 3338) && (pixel_index <= 3339)) || ((pixel_index >= 3347) && (pixel_index <= 3372)) || ((pixel_index >= 3376) && (pixel_index <= 3379)) || ((pixel_index >= 3391) && (pixel_index <= 3397)) || ((pixel_index >= 3403) && (pixel_index <= 3405)) || ((pixel_index >= 3408) && (pixel_index <= 3410)) || pixel_index == 3413 || ((pixel_index >= 3416) && (pixel_index <= 3419)) || pixel_index == 3423 || ((pixel_index >= 3434) && (pixel_index <= 3435)) || pixel_index == 3438 || ((pixel_index >= 3443) && (pixel_index <= 3468)) || ((pixel_index >= 3472) && (pixel_index <= 3475)) || pixel_index == 3484 || ((pixel_index >= 3488) && (pixel_index <= 3490)) || ((pixel_index >= 3492) && (pixel_index <= 3493)) || pixel_index == 3496 || ((pixel_index >= 3500) && (pixel_index <= 3501)) || ((pixel_index >= 3504) && (pixel_index <= 3505)) || pixel_index == 3509 || ((pixel_index >= 3513) && (pixel_index <= 3515)) || ((pixel_index >= 3518) && (pixel_index <= 3520)) || ((pixel_index >= 3524) && (pixel_index <= 3525)) || ((pixel_index >= 3529) && (pixel_index <= 3531)) || ((pixel_index >= 3534) && (pixel_index <= 3535)) || ((pixel_index >= 3539) && (pixel_index <= 3564)) || pixel_index == 3572 || ((pixel_index >= 3580) && (pixel_index <= 3581)) || ((pixel_index >= 3588) && (pixel_index <= 3589)) || ((pixel_index >= 3592) && (pixel_index <= 3593)) || ((pixel_index >= 3596) && (pixel_index <= 3597)) || ((pixel_index >= 3604) && (pixel_index <= 3606)) || ((pixel_index >= 3614) && (pixel_index <= 3616)) || ((pixel_index >= 3620) && (pixel_index <= 3621)) || ((pixel_index >= 3625) && (pixel_index <= 3627)) || ((pixel_index >= 3630) && (pixel_index <= 3631)) || ((pixel_index >= 3635) && (pixel_index <= 3660)) || ((pixel_index >= 3668) && (pixel_index <= 3669)) || ((pixel_index >= 3675) && (pixel_index <= 3678)) || ((pixel_index >= 3683) && (pixel_index <= 3685)) || ((pixel_index >= 3688) && (pixel_index <= 3689)) || pixel_index == 3693 || ((pixel_index >= 3698) && (pixel_index <= 3704)) || ((pixel_index >= 3708) && (pixel_index <= 3712)) || ((pixel_index >= 3715) && (pixel_index <= 3717)) || ((pixel_index >= 3720) && (pixel_index <= 3723)) || ((pixel_index >= 3726) && (pixel_index <= 3728)) || (pixel_index >= 3731) && (pixel_index <= 6143)) oled_data = 16'b1010000000000000;
else if (pixel_index == 2443 || pixel_index == 2449 || pixel_index == 2457 || pixel_index == 2817 || pixel_index == 2834 || pixel_index == 2836 || pixel_index == 3384 || pixel_index == 3426 || pixel_index == 3480 || pixel_index == 3679) oled_data = 16'b1010010100010100;
else if (((pixel_index >= 2447) && (pixel_index <= 2448)) || pixel_index == 2458 || pixel_index == 2530 || pixel_index == 2550 || pixel_index == 2625 || pixel_index == 2749 || pixel_index == 2832 || pixel_index == 2844 || pixel_index == 2989 || pixel_index == 3007 || pixel_index == 3085 || pixel_index == 3181 || pixel_index == 3203 || pixel_index == 3208 || pixel_index == 3222 || pixel_index == 3277 || pixel_index == 3373 || pixel_index == 3469 || pixel_index == 3565 || pixel_index == 3571 || pixel_index == 3661 || pixel_index == 3667) oled_data = 16'b1010001010001010;
else if (pixel_index == 2455) oled_data = 16'b1010001010000000;
else if (pixel_index == 2531 || pixel_index == 2633 || pixel_index == 2635 || pixel_index == 2745 || pixel_index == 2821 || pixel_index == 2828 || pixel_index == 2842 || pixel_index == 3102 || pixel_index == 3324 || pixel_index == 3420 || pixel_index == 3429 || pixel_index == 3508 || pixel_index == 3613 || pixel_index == 3682 || pixel_index == 3697) oled_data = 16'b1010011110011110;
else if (pixel_index == 2538 || pixel_index == 2540 || pixel_index == 2542 || pixel_index == 2544 || ((pixel_index >= 2548) && (pixel_index <= 2549)) || pixel_index == 2552 || pixel_index == 2555 || ((pixel_index >= 2615) && (pixel_index <= 2616)) || pixel_index == 2626 || ((pixel_index >= 2628) && (pixel_index <= 2630)) || pixel_index == 2632 || pixel_index == 2638 || pixel_index == 2640 || pixel_index == 2642 || pixel_index == 2644 || pixel_index == 2646 || pixel_index == 2648 || ((pixel_index >= 2652) && (pixel_index <= 2653)) || ((pixel_index >= 2710) && (pixel_index <= 2714)) || pixel_index == 2722 || ((pixel_index >= 2725) && (pixel_index <= 2726)) || pixel_index == 2728 || pixel_index == 2731 || pixel_index == 2734 || pixel_index == 2736 || pixel_index == 2738 || ((pixel_index >= 2740) && (pixel_index <= 2742)) || pixel_index == 2744 || ((pixel_index >= 2747) && (pixel_index <= 2748)) || pixel_index == 2805 || pixel_index == 2810 || ((pixel_index >= 2818) && (pixel_index <= 2820)) || ((pixel_index >= 2822) && (pixel_index <= 2825)) || pixel_index == 2835 || ((pixel_index >= 2837) && (pixel_index <= 2841)) || pixel_index == 2901 || pixel_index == 2906 || ((pixel_index >= 2990) && (pixel_index <= 2991)) || pixel_index == 2997 || ((pixel_index >= 2999) && (pixel_index <= 3002)) || ((pixel_index >= 3008) && (pixel_index <= 3010)) || ((pixel_index >= 3014) && (pixel_index <= 3015)) || ((pixel_index >= 3018) && (pixel_index <= 3020)) || ((pixel_index >= 3022) && (pixel_index <= 3025)) || ((pixel_index >= 3033) && (pixel_index <= 3035)) || ((pixel_index >= 3039) && (pixel_index <= 3040)) || ((pixel_index >= 3044) && (pixel_index <= 3045)) || ((pixel_index >= 3049) && (pixel_index <= 3050)) || ((pixel_index >= 3052) && (pixel_index <= 3053)) || ((pixel_index >= 3057) && (pixel_index <= 3058)) || ((pixel_index >= 3086) && (pixel_index <= 3087)) || ((pixel_index >= 3093) && (pixel_index <= 3098)) || ((pixel_index >= 3103) && (pixel_index <= 3107)) || ((pixel_index >= 3110) && (pixel_index <= 3111)) || ((pixel_index >= 3114) && (pixel_index <= 3115)) || ((pixel_index >= 3118) && (pixel_index <= 3123)) || ((pixel_index >= 3127) && (pixel_index <= 3133)) || ((pixel_index >= 3135) && (pixel_index <= 3136)) || ((pixel_index >= 3140) && (pixel_index <= 3141)) || ((pixel_index >= 3144) && (pixel_index <= 3146)) || ((pixel_index >= 3148) && (pixel_index <= 3150)) || ((pixel_index >= 3153) && (pixel_index <= 3154)) || ((pixel_index >= 3182) && (pixel_index <= 3183)) || ((pixel_index >= 3188) && (pixel_index <= 3195)) || ((pixel_index >= 3197) && (pixel_index <= 3199)) || ((pixel_index >= 3206) && (pixel_index <= 3207)) || ((pixel_index >= 3209) && (pixel_index <= 3210)) || ((pixel_index >= 3214) && (pixel_index <= 3215)) || ((pixel_index >= 3218) && (pixel_index <= 3220)) || ((pixel_index >= 3223) && (pixel_index <= 3224)) || ((pixel_index >= 3228) && (pixel_index <= 3229)) || ((pixel_index >= 3232) && (pixel_index <= 3233)) || ((pixel_index >= 3235) && (pixel_index <= 3238)) || ((pixel_index >= 3240) && (pixel_index <= 3241)) || ((pixel_index >= 3244) && (pixel_index <= 3247)) || ((pixel_index >= 3249) && (pixel_index <= 3250)) || ((pixel_index >= 3278) && (pixel_index <= 3279)) || ((pixel_index >= 3284) && (pixel_index <= 3287)) || ((pixel_index >= 3289) && (pixel_index <= 3291)) || ((pixel_index >= 3293) && (pixel_index <= 3294)) || ((pixel_index >= 3302) && (pixel_index <= 3305)) || ((pixel_index >= 3310) && (pixel_index <= 3311)) || ((pixel_index >= 3315) && (pixel_index <= 3316)) || ((pixel_index >= 3318) && (pixel_index <= 3319)) || ((pixel_index >= 3325) && (pixel_index <= 3326)) || ((pixel_index >= 3328) && (pixel_index <= 3329)) || ((pixel_index >= 3331) && (pixel_index <= 3334)) || ((pixel_index >= 3336) && (pixel_index <= 3337)) || ((pixel_index >= 3340) && (pixel_index <= 3346)) || ((pixel_index >= 3374) && (pixel_index <= 3375)) || ((pixel_index >= 3380) && (pixel_index <= 3383)) || ((pixel_index >= 3385) && (pixel_index <= 3387)) || ((pixel_index >= 3389) && (pixel_index <= 3390)) || ((pixel_index >= 3398) && (pixel_index <= 3402)) || ((pixel_index >= 3406) && (pixel_index <= 3407)) || ((pixel_index >= 3411) && (pixel_index <= 3412)) || ((pixel_index >= 3414) && (pixel_index <= 3415)) || ((pixel_index >= 3421) && (pixel_index <= 3422)) || ((pixel_index >= 3424) && (pixel_index <= 3425)) || pixel_index == 3427 || pixel_index == 3430 || pixel_index == 3432 || ((pixel_index >= 3436) && (pixel_index <= 3437)) || ((pixel_index >= 3439) && (pixel_index <= 3442)) || ((pixel_index >= 3470) && (pixel_index <= 3471)) || ((pixel_index >= 3476) && (pixel_index <= 3479)) || ((pixel_index >= 3481) && (pixel_index <= 3483)) || ((pixel_index >= 3485) && (pixel_index <= 3487)) || ((pixel_index >= 3494) && (pixel_index <= 3495)) || ((pixel_index >= 3497) && (pixel_index <= 3498)) || ((pixel_index >= 3502) && (pixel_index <= 3503)) || ((pixel_index >= 3506) && (pixel_index <= 3507)) || ((pixel_index >= 3511) && (pixel_index <= 3512)) || ((pixel_index >= 3516) && (pixel_index <= 3517)) || ((pixel_index >= 3521) && (pixel_index <= 3523)) || ((pixel_index >= 3526) && (pixel_index <= 3528)) || ((pixel_index >= 3532) && (pixel_index <= 3533)) || ((pixel_index >= 3536) && (pixel_index <= 3538)) || ((pixel_index >= 3566) && (pixel_index <= 3570)) || ((pixel_index >= 3573) && (pixel_index <= 3579)) || ((pixel_index >= 3582) && (pixel_index <= 3587)) || ((pixel_index >= 3590) && (pixel_index <= 3591)) || ((pixel_index >= 3594) && (pixel_index <= 3595)) || ((pixel_index >= 3598) && (pixel_index <= 3603)) || ((pixel_index >= 3607) && (pixel_index <= 3612)) || ((pixel_index >= 3617) && (pixel_index <= 3619)) || ((pixel_index >= 3622) && (pixel_index <= 3624)) || ((pixel_index >= 3628) && (pixel_index <= 3629)) || ((pixel_index >= 3633) && (pixel_index <= 3634)) || ((pixel_index >= 3662) && (pixel_index <= 3666)) || ((pixel_index >= 3670) && (pixel_index <= 3674)) || ((pixel_index >= 3680) && (pixel_index <= 3681)) || ((pixel_index >= 3686) && (pixel_index <= 3687)) || ((pixel_index >= 3691) && (pixel_index <= 3692)) || ((pixel_index >= 3694) && (pixel_index <= 3696)) || ((pixel_index >= 3705) && (pixel_index <= 3707)) || ((pixel_index >= 3713) && (pixel_index <= 3714)) || ((pixel_index >= 3718) && (pixel_index <= 3719)) || ((pixel_index >= 3724) && (pixel_index <= 3725)) || (pixel_index >= 3729) && (pixel_index <= 3730)) oled_data = 16'b1111011110011110;
else if (pixel_index == 2547 || pixel_index == 2557 || pixel_index == 2709 || pixel_index == 2730) oled_data = 16'b0101000000000000;
else if (pixel_index == 2556 || pixel_index == 2733 || pixel_index == 2827 || pixel_index == 2907 || pixel_index == 2998 || pixel_index == 3003 || pixel_index == 3099 || pixel_index == 3113 || pixel_index == 3288 || pixel_index == 3431 || pixel_index == 3491 || pixel_index == 3499) oled_data = 16'b1111011110010100;
else if (pixel_index == 2636 || pixel_index == 2746) oled_data = 16'b1111010100011110;
else if (pixel_index == 2645 || pixel_index == 2650 || pixel_index == 2724 || pixel_index == 2729 || pixel_index == 2826 || pixel_index == 2843 || pixel_index == 3428 || pixel_index == 3433 || pixel_index == 3510 || pixel_index == 3632) oled_data = 16'b1111010100010100;
else if (pixel_index == 3388) oled_data = 16'b1010010100001010;
else if (pixel_index == 3690) oled_data = 16'b1010011110010100;
else oled_data = 0;
end
    
endmodule
