`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 22.03.2022 00:31:03
// Design Name: 
// Module Name: menu
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module menu(input pbu, pbd, SW0, input [31:0] x, y, input clk, input [3:0] layer, output reg [15:0] oled_data, output reg [3:0] state);
    parameter [31:0]a = 3;
    parameter [31:0]b = 12;
    parameter [31:0]c = 12;
    parameter [31:0]d = 22;
    parameter [31:0]e = 29;
    parameter [31:0]f = 39;
    wire [15:0] menudisp [5:0];
    wire vert, vert2, vert3, welcome, trace, distance, arrow1, arrow2, arrow3, arrow4, landmarks, labtask, timer;
    wire boxwidth, box1, box2, box3, box4, box5;

    assign vert = y >= 25 && y <= 31;
    assign vert2 = y >= 39 && y <= 45;
    assign vert3 = y >= 53 && y <= 59;
    assign welcome = (y == a && (x == 29 ||  x == 33 || (x >= 35 && x <= 39) || x == 41 || (x >= 48 && x <= 50) || (x >= 54 && x <= 56) || x == 59 || x == 63 || (x >= 65 && x <= 69) || x == 72))
              || (y == a + 1 && (x == 29 ||  x == 33 || x == 35 || x == 41 || x == 47 || x == 51 || x == 53 || x == 57 || x == 59 || x == 60 || x == 62 || x == 63 || x == 65 || x == 72))
              || (y == a + 2 && (x == 29 ||  x == 33 || x == 35 || x == 41 || x == 47 || x == 53 || x == 57 || x == 59 || x == 61 || x == 63 || x == 65 || x == 72))
              || (y == a + 3 && (x == 29 ||  x == 33 || (x >= 35 && x <= 37) || x == 41 || x == 47 || x == 53 || x == 57 || x == 59 || x == 63 || (x >= 65 && x <= 67) || x == 72))
              || (y == a + 4 && (x == 29 ||  x == 31 ||  x == 33 || x == 35 || x == 41 || x == 47 || x == 53 || x == 57 || x == 59 || x == 63 || x == 65 || x == 72))
              || (y == a + 5 && (x == 29 ||  x == 31 ||  x == 33 || x == 35 || x == 41 || x == 47 || x == 51 || x == 53 || x == 57 || x == 59 || x == 63 || x == 65))
              || (y == a + 6 && (x == 30 ||  x == 32 || (x >= 35 && x <= 39) || (x >= 41 && x <= 45) || (x >= 48 && x <= 50) || (x >= 54 && x <= 56) || x == 57 || x == 59 || x == 63 || (x >= 65 && x <= 69) || x == 72))
              || (y == a + 10 && ((x >= 16 && x <= 19) || x == 22 || (x >= 25 && x <= 27) || x == 30 || x == 34 || x == 40 || x == 44 || x == 48 || (x >= 53 && x <= 55) || (x >= 58 && x <= 61) || (x >= 64 && x <= 68) || x == 70 || (x >= 73 && x <= 75) || x == 78 || x == 82 || x == 84))
              || (y == a + 11 && (x == 16 || x == 20 || x == 22 || x == 24 || x == 28 || x == 30 || x == 34 || x == 39 || x == 41 || x == 44 || x == 48 || x == 52 || x == 56 || x == 58 || x == 62 || x == 66 || x == 70 || x == 72 || x == 76 || x == 78 || x == 82 || x == 84))
              || (y == a + 12 && (x == 16 || x == 20 || x == 22 || x == 24 || x == 30 || x == 33 || x == 38 || x == 42 || x == 44 || x == 45 || x == 48 || x == 52 || x == 56 || x == 58 || x == 62 || x == 66 || x == 70 || x == 72 || x == 76 || x == 78 || x == 79 || x == 82 || x == 84)) 
              || (y == a + 13 && ((x >= 16 && x <= 19) || x == 22 || x == 24 || (x >= 30 && x <= 32) || x == 38 || x == 42 || x == 44 || x == 46 || x == 48 || x == 52 || x == 56 || (x >= 58 && x <= 61) || x == 66 || x == 70 || x == 72 || x == 76 || x == 78 || x == 80 || x == 82 || x == 84))
              || (y == a + 14 && (x == 16 || x == 22 || x == 24 || x == 30 || x == 33 || (x >= 38 && x <= 42) || x == 44 || x == 47 || x == 48 || x == 52 || x == 56 || x == 58 || x == 66 || x == 70 || x == 72 || x == 76 || x == 78 || x == 81 || x == 82 || x == 84)) 
              || (y == a + 15 && (x == 16 || x == 22 || x == 24 || x == 28 || x == 30 || x == 34 || x == 38 || x == 42 || x == 44 || x == 48 || x == 52 || x == 56 || x == 58 || x == 66 || x == 70 || x == 72 || x == 76 || x == 78 || x == 82))
              || (y == a + 16 && (x == 16 || x == 22 || (x >= 25 && x <= 27) || x == 30 || x == 34 || x == 38 || x == 42 || x == 44 || x == 48 || (x >= 53 && x <= 55) || x == 58 || x == 66 || x == 70 || (x >= 73 && x <= 75) || x == 78 || x == 82 || x == 84));

    assign distance = (x == b && (y >= 25 && y <= 31)) || (x == b + 1 && (y == 25 || y == 31)) || (x == b + 2 && (y == 25 || y == 31)) || (x == b + 2 && (y == 25 || y == 31)) || (x == b + 3 && (y == 25 || y == 31)) || (x == b + 4 && (y >= 26 && y <= 30))
             || (x == b + 6 && (y >= 25 && y <= 31))
             || (x == b + 8 && (y == 26 || y == 27 || y == 30)) || (x == b + 9 && (y == 25 || y == 28 || y == 31)) || (x == b + 10 && (y == 25 || y == 28 || y == 31)) || (x == b + 11 && (y == 25 || y == 28 || y == 31)) || (x == b + 12 && (y == 26 || y == 29 || y == 30)) 
             || (x == b + 14 && y == 25) || (x == b + 15 && y == 25) || (x == b + 16 && (y >= 25 && y <= 31)) || (x == b + 17 && y == 25) || (x == b + 18 && y == 25)
             || (x == b + 20 && (y >= 27 && y <= 31)) || (x == b + 21 && (y == 26 || y == 29)) || (x == b + 22 && (y == 25 || y == 29)) || (x == b + 23 && (y == 26 || y == 29)) || (x == b + 24 && (y >= 27 && y <= 31))
             || (x == b + 26 && (y >= 25 && y <= 31)) || (x == b + 27 && y == 26) || (x == b + 28 && y == 27) || (x == b + 29 && y == 28) || (x == b + 30 && (y >= 25 && y <= 31))
             || (x == b + 32 && (y >= 26 && y <= 30)) || (x == b + 33 && (y == 25 || y == 31)) || (x == b + 34 && (y == 25 || y == 31)) || (x == b + 35 && (y == 25 || y == 31)) || (x == b + 36 && (y == 26 || y == 30))
             || (x == b + 38 && (y >= 25 && y <= 31)) || (x == b + 39 && (y == 25 || y == 28 || y == 31)) || (x == b + 40 && (y == 25 || y == 28 || y == 31)) || (x == b + 41 && (y == 25 || y == 31)) || (x == b + 42 && (y == 25 || y == 31))
             || (x == b + 48 && vert) || (x == b + 49 && (y == 25 || y == 28)) || (x == b + 50 && (y == 25 || y == 28)) || (x == b + 51 && y == 25) || (x == b + 52 && y == 25)
             || (x == b + 54 && (y >= 25 && y <= 31))
             || (x == b + 56 && (y >= 25 && y <= 31)) || (x == b + 57 && y == 26) || (x == b + 58 && y == 27) || (x == b + 59 && y == 28) || (x == b + 60 && (y >= 25 && y <= 31))
             || (x == b + 62 && (y >= 25 && y <= 31)) || (x == b + 63 && (y == 25 || y == 31)) || (x == b + 64 && (y == 25 || y == 31)) || (x == b + 65 && (y == 25 || y == 31)) || (x == b + 66 && (y == 25 || y == 31)) || (x == b + 67 && (y >= 26 && y <= 30))
             || (x == b + 69 && (y >= 25 && y <= 31)) || (x == b + 70 && (y == 25 || y == 28 || y == 31)) || (x == b + 71 && (y == 25 || y == 28 || y == 31)) || (x == b + 72 && (y == 25 || y == 31)) || (x == b + 73 && (y == 25 || y == 31))
             || (x == b + 75 && vert) || (x == b + 76 && (y == 25 || y == 28)) || (x == b + 77 && (y == 25 || y == 28 || y == 29)) || (x == b + 78 && (y == 25 || y == 28 || y == 30)) || (x == b + 79 && (y == 26 || y == 27 || y == 31));
             
     assign trace = (x == c && y == 39) || (x == c + 1 && y == 39) || (x == c + 2 && (y >= 39 && y <= 45)) || (x == c + 3 && y == 39) || (x == c + 4 && y == 39)
                  || (x == c + 6 && vert2) || (x == c + 7 && (y == 39 || y == 42)) || (x == c + 8 && (y == 39 || y == 42 || y == 43)) || (x == c + 9 && (y == 39 || y == 42 || y == 44)) || (x == c + 10 && (y == 40 || y == 41 || y == 45))
                  || (x == c + 12 && (y >= 41 && y <= 45)) || (x == c + 13 && (y == 40 || y == 43)) || (x == c + 14 && (y == 39 || y == 43)) || (x == c + 15 && (y == 40 || y == 43)) || (x == c + 16 && (y >= 41 && y <= 45))
                  || (x == c + 18 && (y >= 40 && y <= 44)) || (x == c + 19 && (y == 39 || y == 45)) || (x == c + 20 && (y == 39 || y == 45)) || (x == c + 21 && (y == 39 || y == 45)) || (x == c + 22 && (y == 40 || y == 44))
                  || (x == c + 24 && vert2) || (x == c + 25 && (y == 39 || y == 42 || y == 45)) || (x == c + 26 && (y == 39 || y == 42 || y == 45)) || (x == c + 27 && (y == 39 || y == 45)) || (x == c + 28 && (y == 39 || y == 45))
                  || (x == c + 32 && y == 39) || (x == c + 33 && y == 39) || (x == c + 34 && (y >= 39 && y <= 45)) || (x == c + 35 && y == 39) || (x == c + 36 && y == 39)
                  || (x == c + 38 && (y >= 40 && y <= 44)) || (x == c + 39 && (y == 39 || y == 45)) || (x == c + 40 && (y == 39 || y == 45)) || (x == c + 41 && (y == 39 || y == 45)) || (x == c + 42 && (y >= 40 && y <= 44))
                  || (x == c + 44 && (y >= 40 && y <= 44)) || (x == c + 45 && (y == 39 || y == 45)) || (x == c + 46 && (y == 39 || y == 42 || y == 45)) || (x == c + 47 && (y == 39 || y == 42 || y == 45)) || (x == c + 48 && (y == 40 || y == 43 || y == 44))
                  || (x == c + 50 && (y >= 39 && y <= 45)) || (x == c + 51 && (y == 39 || y == 42 || y == 45)) || (x == c + 52 && (y == 39 || y == 42 || y == 45)) || (x == c + 53 && (y == 39 || y == 45)) || (x == c + 54 && (y == 39 || y == 45))
                  || (x == c + 56 && y == 39) || (x == c + 57 && y == 39) || (x == c + 58 && (y >= 39 && y <= 45)) || (x == c + 59 && y == 39) || (x == c + 60 && y == 39)
                  || (x == c + 62 && vert2) || (x == c + 63 && y == 42) || (x == c + 64 && y == 42) || (x == c + 65 && y == 42) || (x == c + 66 && vert2)
                  || (x == c + 68 && (y >= 39 && y <= 45)) || (x == c + 69 && (y == 39 || y == 42 || y == 45)) || (x == c + 70 && (y == 39 || y == 42 || y == 45)) || (x == c + 71 && (y == 39 || y == 45)) || (x == c + 72 && (y == 39 || y == 45))
                  || (x == c + 74 && vert2) || (x == c + 75 && (y == 39 || y == 42)) || (x == c + 76 && (y == 39 || y == 42 || y == 43)) || (x == c + 77 && (y == 39 || y == 42 || y == 44)) || (x == c + 78 && (y == 40 || y == 41 || y == 45));
 
    assign landmarks = (x == d && vert3) || (x == d+1 && y == 59) || (x == d+2 && y == 59) || (x == d+3 && y == 59) || (x == d+4 && y == 59) 
    || (x == d+6 && (y >= 55 && y <= 59)) || (x == d+7 && (y == 54 || y == 57)) || (x == d+8 && (y == 53 || y == 57)) || (x == d+9 && (y == 54 || y == 57)) || (x == d+10 && (y >= 55 && y <= 59))
    || (x == d+12 && vert3) || (x == d+13 && y == 55) || (x == d+14 && y == 56) || (x == d+15 && y == 57) || (x == d+16 && vert3)
    || (x == d+18 && vert3) || (x == d+19 && (y == 53 || y == 59)) || (x == d+20 && (y == 53 || y == 59)) || (x == d+21 && (y == 53 || y == 59)) || (x == d+22 && (y >= 54 && y <= 58))
    || (x == d+24 && vert3) || (x == d+25 && y == 54) || (x == d+26 && y == 55) || (x == d+27 && y == 54) || (x == d+28 && vert3)
    || (x == d+30 && (y >= 55 && y <= 59)) || (x == d+31 && (y == 54 || y == 57)) || (x == d+32 && (y == 53 || y == 57)) || (x == d+33 && (y == 54 || y == 57)) || (x == d+34 && (y >= 55 && y <= 59))
    || (x == d+36 && vert3) || (x == d+37 && (y == 53 || y == 56)) || (x == d+38 && (y == 53 || y == 56 || y == 57)) || (x == d+39 && (y == 53 || y == 56 || y == 58)) || (x == d+40 && (y == 54 || y == 55 || y == 59))
    || (x == d+42 && vert3) || (x == d+43 && y == 56) || (x == d+44 && y == 56) || (x == d+45 && (y == 55 || y == 57)) || (x == d+46 && (y == 53 || y == 54 || y == 58 || y == 59))
    || (x == d+48 && (y == 54 || y == 55 || y == 58)) || (x == d+49 && (y == 53 || y == 56 || y == 59)) || (x == d+50 && (y == 53 || y == 56 || y == 59)) || (x == d+51 && (y == 53 || y == 56 || y == 59)) || (x == d+52 && (y == 54 || y == 57 || y == 58));
    
    assign labtask = (x == e && (y >= 25 && y <= 31)) || (x==e+1 && y==31) || (x==e+2 && y==31) || (x==e+3 && y==31) || (x==e+4 && y==31)
                    || (x == e + 6 && (y >= 27 && y <= 31)) || (x == e + 7 && (y == 26 || y == 29)) || (x == e + 8 && (y == 25 || y == 29)) || (x == e + 9 && (y == 26 || y == 29)) || (x == e + 10 && (y >= 27 && y <= 31))
                    || (x == e+12 && (y >= 25 && y <= 31)) || (x == e+13 && (y == 25 || y==28 || y == 31)) || (x == e+14 && (y == 25 || y==28 || y == 31)) || (x == e+15 && (y == 25 || y==28 || y == 31)) || (x == e+16 && (y == 26 || y==27 || y==29 || y == 30))
                    || (x == e + 21 && y == 25) || (x == e + 22 && y == 25) || (x == e + 23 && (y >= 25 && y <= 31)) || (x == e + 24 && y == 25) || (x == e + 25 && y == 25)
                    || (x == e + 27 && (y >= 27 && y <= 31)) || (x == e + 28 && (y == 26 || y == 29)) || (x == e + 29 && (y == 25 || y == 29)) || (x == e + 30 && (y == 26 || y == 29)) || (x == e + 31 && (y >= 27 && y <= 31))
                    || (x == e + 33 && (y == 26 || y == 27 || y == 30)) || (x == e + 34 && (y == 25 || y == 28 || y == 31)) || (x == e + 35 && (y == 25 || y == 28 || y == 31)) || (x == e + 36 && (y == 25 || y == 28 || y == 31)) || (x == e + 37 && (y == 26 || y == 29 || y == 30)) 
                    || (x == e+39 && vert) || (x==e+40 && y==28) || (x==e+41 && y==28) || (x==e+42 && (y==27 || y==29)) || (x==e+43 && (y==25 || y==30 || y==26 || y==31));
     
     assign timer =  (x == f && y == 39) || (x == f + 1 && y == 39) || (x == f + 2 && (y >= 39 && y <= 45)) || (x == f + 3 && y == 39) || (x == f + 4 && y == 39)
                    || (x == f + 6 && vert2) 
                    || (x == f + 8 && vert2) || (x == f + 9 && y==40) || (x == f + 10 && y==41) || (x == f + 11 && y==40) || (x == f + 12 && vert2)
                    || (x == f + 14 && vert2) || (x == f + 15 && (y == 39 || y == 42 || y == 45)) || (x == f + 16 && (y == 39 || y == 42 || y == 45)) || (x == f + 17 && (y == 39 || y == 45)) || (x == f + 18 && (y == 39 || y == 45))
                    || (x == f + 20 && vert2) || (x == f + 21 && (y == 39 || y == 42)) || (x == f + 22 && (y == 39 || y == 42 || y == 43)) || (x == f + 23 && (y == 39 || y == 42 || y == 44)) || (x == f + 24 && (y == 40 || y == 41 || y == 45));

              
    
    assign boxwidth = (x >= 0 && x <= 95);
    assign arrow1 = (((y >= 25 && y <= 31) && x == 4) || (x == 5 && (y == 25 || y == 31))  || (x == 6 && (y == 26 || y == 30)) || (x == 7 && (y == 27 || y == 29)) || x == 8 && y == 28);
    assign arrow2 = (((y >= 39 && y <= 45) && x == 4) || (x == 5 && (y == 39 || y == 45))  || (x == 6 && (y == 40 || y == 44)) || (x == 7 && (y == 41 || y == 43)) || x == 8 && y == 42);
    assign arrow3 = (((y >= 53 && y <= 59) && x == 4) || (x == 5 && (y == 53 || y == 59))  || (x == 6 && (y == 54 || y == 58)) || (x == 7 && (y == 55 || y == 57)) || x == 8 && y == 56);
    
    assign box1 = ((y >= 23 && y <= 33) && boxwidth && ~distance && ~arrow1);
    assign box2 = ((y >= 37 && y <= 47) && boxwidth && ~trace && ~arrow2);
    assign box3 = ((y >= 51 && y <= 61) && boxwidth && ~landmarks && ~arrow3);
    assign box4 = ((y >= 23 && y <= 33) && boxwidth && ~labtask && ~arrow1);
    assign box5 = ((y >= 37 && y <= 47) && boxwidth && ~timer && ~arrow2);
    
    assign menudisp[0] = (welcome || distance || trace || landmarks);
    assign menudisp[1] = (welcome || trace || landmarks || box1);
    assign menudisp[2] = (welcome || distance || landmarks || box2);
    assign menudisp[3] = (welcome || distance || trace || box3);
    assign menudisp[4] = (welcome || box4 || timer);
    assign menudisp[5] = (welcome || box5 || labtask);
    
    always @ (posedge clk) begin
        state <= pbu && layer == 0 && state != 0 ? state - 1 : pbd && layer == 0 && state != 5 ? state + 1 : state;
    end
    
    always @ (*) begin
        if(SW0 && layer == 0)
           oled_data = menudisp[state] ? 16'b1111100000000000 : 16'b1111111111111111;
        else
           oled_data = menudisp[state] ? 16'b1111111111111111 : 16'b1111100000000000; 
    end 
    
endmodule
